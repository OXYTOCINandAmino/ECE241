
module Divider(SW, KEY, CLOCK_50,HEX0, HEX2,HEX4,HEX5);
    input [7:0] SW;
    input [1:0] KEY;
    input CLOCK_50;
   
    output [6:0] HEX0, HEX2,HEX4,HEX5;

    wire reset;
    wire go;
	 
	 wire [3:0]Divisor;
	 wire [3:0]divident;
	 wire [3:0]Quotient;
	 wire [3:0]Remainder;

    assign go = ~KEY[1];
    assign reset = KEY[0];
	 assign clk=CLOCK_50;

    part3 u0(
        .clk(clk),
        .reset(reset),
        .go(go),
        .Divisor(Divisor),
	     .divident(divident),
	     .Quotient(Quotient),
	     .Remainder(Remainder)
    );
      
 

    hex_decoder H0(
        .hex_digit(Divisor), 
        .segments(HEX0)
        );
        
    hex_decoder H1(
        .hex_digit(divident), 
        .segments(HEX2)
        );
    hex_decoder H2(
        .hex_digit(Quotient), 
        .segments(HEX4)
        );
        
    hex_decoder H3(
        .hex_digit(Remainder), 
        .segments(HEX5)
        );	

endmodule


module part3(
    input clk,
    input reset,
    input go,
    input [3:0]Divisor,
	 input [3:0]divident,
	 output [3:0]Quotient,
	 output [3:0]Remainder
    );
//
wire ld;
wire ld_final;
wire Shift_L;
wire Subtract;
wire [4:0]remainder;
assign Remainder[3:0]=remainder[3:0];
    

    control C0(
    .clk(clk),
    .reset(reset),
    .go(go),
    .ld(ld),
	 .ld_final(ld_final),
    .Shift_L(Shift_L),
	 .Subtract(Subtract)
    );
	 //

    datapath D0(
	 .clk(clk),
	 .reset(reset),
	 .ld(ld),
	 .ld_final(ld_final),
    .Divisor(Divisor),
	 .divident(divident),
    .Shift_L(Shift_L),
	 .Subtract(Subtract),
	 .Reg_A_Final(remainder),
	 .Divident_Final(Quotient)
	 );
                
 endmodule 
////////////////////////////////////////////////////////////////
module control(
    input clk,
    input reset,
    input go,

    output reg  ld,ld_final,
    output reg  Shift_L,Subtract
    );

    reg [5:0] current_state, next_state; 
    
    localparam  S_LOAD        = 5'd0,
                S_LOAD_WAIT   = 5'd1,
					 
					 Operate_1 = 5'd2,
					 Load_Back_1 = 5'd3,
					 
					 Operate_2 = 5'd4,
					 Load_Back_2 = 5'd5,
					 
					 Operate_3 = 5'd6,
					 Load_Back_3 = 5'd7,
					 
					 Operate_Final = 5'd8;
   
    
    // Next state logic aka our state table
	
    always@(*)
    begin: state_table 
            case (current_state)
                S_LOAD: next_state = go ? S_LOAD_WAIT : S_LOAD; // Loop in current state until value is input
                S_LOAD_WAIT: next_state = go ? S_LOAD_WAIT : Operate_1 ; // Loop in current state until go signal goes low
                
					 Operate_1:   next_state = Load_Back_1;
					 Load_Back_1: next_state = Operate_2;
					 Operate_2:   next_state = Load_Back_2;
					 Load_Back_2: next_state = Operate_3;
					 Operate_3:   next_state = Load_Back_3;
					 Load_Back_3: next_state = Operate_Final;
			   Operate_Final:   next_state = S_LOAD;
                // we will be done our two operations, start over after
            default:     next_state = S_LOAD;
        endcase
    end
 //
 
    always @(*)
    begin: enable_signals
        // By default make all our signals 0 to avoid latches.
        // This is a different style from using a default statement.
        // It makes the code easier to read.  If you add other out
        // signals be sure to assign a default value for them here.
        ld = 1'b0;
        ld_final = 1'b0;
        Shift_L=1'b 0;
		  Subtract=1'b 0;
		  
        case (current_state)
            S_LOAD: begin
                ld = 1'b1;
                end
		
				Operate_1:
				    begin
					 Shift_L= 1'b1;
					 Subtract = 1'b1;
					 end
				Load_Back_1:
					 begin
					 ld = 1'b1;
					 ld_final=1'b1;
					 end
		      Operate_2:
				    begin
					 Shift_L= 1'b1;
					 Subtract = 1'b1;
					 end
				Load_Back_2:
					 begin
					 ld = 1'b1;
					 ld_final=1'b1;
					 end
			   Operate_3:
				    begin
					 Shift_L= 1'b1;
					 Subtract = 1'b1;
					 end
				Load_Back_3:
					 begin
					 ld = 1'b1;
					 ld_final=1'b1;
					 end
				Operate_Final:
				    begin
					 Shift_L= 1'b1;
					 Subtract = 1'b1;
					 end
					 
        endcase
    end // enable_signals
   
    // current_state registers
    always@(posedge clk)
    begin: state_FFs
        if(reset)
            current_state <= S_LOAD;
        else
            current_state <= next_state;
    end // state_FFS
endmodule
					 

///////////////////////////////////////////////////////////////
module datapath(clk,reset,ld,ld_final,
                 Divisor,divident,
                 Shift_L,Subtract,
					  Reg_A_Final,Divident_Final);

input clk;
input reset;

input [4:0]Divisor;
input [3:0]divident;

input ld, ld_final;
input Shift_L;
input Subtract;

//output
output reg [4:0]Reg_A_Final;
output reg [3:0]Divident_Final;

//registers
reg [4:0]Reg_A;
reg [3:0]Divident;
wire  [4:0]reg_A= 5'b 0;
   
always@(posedge clk) begin
        if(reset==1) begin
             Reg_A <= 5'b 0;
		       Divident <= 4'b 0;
        end
        else begin
            if(ld==1)
	         Reg_A <= ld_final ? Reg_A_Final : reg_A;
		      Divident <= ld_final ? Divident_Final : divident;
        end
    end	
//shift Left
reg [4:0]Reg_A_shift;
reg [3:0]Divident_shift;

always @(*)
	begin
	if(Shift_L==1)
	   begin
	   Reg_A_shift = Reg_A<<1;
		Reg_A_shift[0] = Divident[3];
		Divident_shift = Divident<<1;
		end
	end
//


	//Subtract
reg [4:0]Reg_A_subtract;
always @(*)
	begin
	if(Subtract==1)
	   begin
	   Reg_A_subtract = Reg_A_shift - Divisor;
		end
	end
//

//Reg_A Divident Final 


always @(*)
	begin
	if(Reg_A_subtract[4]==1)
	   begin
	   Reg_A_Final = Reg_A_shift;
		Divident_Final= Divident_shift;
		end
		
	else if(Reg_A_subtract[4]==0)
	   begin
	   Reg_A_Final = Reg_A_subtract;
		Divident_Final= Divident_shift;
		Divident_Final[0]=1;
		end
	end
//


endmodule

module hex_decoder(hex_digit, segments);
    input [3:0] hex_digit;
    output reg [6:0] segments;
   
    always @(*)
        case (hex_digit)
            4'h0: segments = 7'b100_0000;
            4'h1: segments = 7'b111_1001;
            4'h2: segments = 7'b010_0100;
            4'h3: segments = 7'b011_0000;
            4'h4: segments = 7'b001_1001;
            4'h5: segments = 7'b001_0010;
            4'h6: segments = 7'b000_0010;
            4'h7: segments = 7'b111_1000;
            4'h8: segments = 7'b000_0000;
            4'h9: segments = 7'b001_1000;
            4'hA: segments = 7'b000_1000;
            4'hB: segments = 7'b000_0011;
            4'hC: segments = 7'b100_0110;
            4'hD: segments = 7'b010_0001;
            4'hE: segments = 7'b000_0110;
            4'hF: segments = 7'b000_1110;   
            default: segments = 7'h7f;
        endcase
endmodule






////////////////////////////////////////////////////////////////
module show_part3(input clk,
    input reset,
    input go,
    input [3:0]Divisor,
	 input [3:0]divident,
	 input [3:0]Quotient,
	 input [3:0]Remainder);
	 wire ld;
    wire ld_final;
    wire Shift_L;
    wire Subtract;
	  control C0(
    .clk(clk),
    .reset(reset),
    .go(go),
    .ld(ld),
	 .ld_final(ld_final),
    .Shift_L(Shift_L),
	 .Subtract(Subtract)
    );
	 endmodule
////////////////////////////////////////////////////////////////