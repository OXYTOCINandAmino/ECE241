module ratedivider(enable, load, clk, reset_n, q);
	input enable, clk, reset_n;
	input [2:0] load;
	output reg [2:0] q;
	
	always @(posedge clk)
	begin
		if (reset_n == 1'b0)
			q <= load;
		else if (enable == 1'b1)
			begin
				if (q == 0)
					q <= load;
				else
					q <= q - 1'b1;
			end
	end
endmodule

